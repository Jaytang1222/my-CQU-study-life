`timescale 1ns / 1ps

module nxor_sim();
    // 输入信号定义
    reg [31:0] a;
    reg [31:0] b;
    
    // 输出信号定义
    wire [31:0] c;
    
    // 实例化32位同或门（使用参数化模块）
    norgate #(.WIDTH(32)) uut (
        .a(a),
        .b(b),
        .c(c)
    );
    
    // 监控信号变化
    initial begin
        $monitor("时间 = %0t, a = %h, b = %h, 输出c = %h", $time, a, b, c);
    end
    
    // 测试序列
    initial begin
        // 初始化输入
        a = 32'h00000000;
        b = 32'h00000000;
        #100;
        
        // 测试1：全0输入（预期输出全1）
        a = 32'h00000000;
        b = 32'h00000000;
        #100;
        
        // 测试2：a全1，b全0（预期输出全0）
        a = 32'hFFFFFFFF;
        b = 32'h00000000;
        #100;
        
        // 测试3：a全0，b全1（预期输出全0）
        a = 32'h00000000;
        b = 32'hFFFFFFFF;
        #100;
        
        // 测试4：全1输入（预期输出全1）
        a = 32'hFFFFFFFF;
        b = 32'hFFFFFFFF;
        #100;
        
        // 测试5：交替位模式（预期输出全0）
        a = 32'hAAAAAAAA;
        b = 32'h55555555;
        #100;
        
        // 测试6：部分位相同模式（预期相同位为1，不同位为0）
        a = 32'h12345678;
        b = 32'h12345678;
        #100;
        
        // 测试7：随机差异模式
        a = 32'h12345678;
        b = 32'h1234ABCD;
        #100;
        
        // 结束仿真
        $finish;
    end
endmodule
